`default_nettype none
/* This is the ps2 port interface for a keyboard.
 *
 */
module key_ctrl();
  
  input clk; // needs to be between 20kHz and 33.3 kHz
  
