// Dummy 